`include "memory.sv"
`include "mem_comm.sv"
`include "mem_tx.sv"
`include "mem_gen.sv"
`include "mem_intrf.sv"
`include "mem_bfm.sv"
`include "mem_mon.sv"
`include "mem_cov.sv"
`include "mem_agent.sv"
`include "mem_sbd.sv"
`include "mem_env.sv"
`include "mem_assert.sv"
`include "mem_tb.sv"
